
module ROM_RS_tx_UE0_real (
	address,
	clock,
	q);	

	input	[10:0]	address;
	input		clock;
	output	[17:0]	q;
endmodule
